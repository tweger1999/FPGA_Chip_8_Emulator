----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 02/25/2023 02:52:56 PM
-- Design Name: 
-- Module Name: FX33 - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity FX33 is
    Port ( Data_In : in STD_LOGIC_VECTOR (7 downto 0);
           X : out STD_LOGIC_VECTOR (7 downto 0);
           Y : out STD_LOGIC_VECTOR (7 downto 0);
           N : out STD_LOGIC_VECTOR (7 downto 0));
end FX33;

architecture Behavioral of FX33 is
begin

process(data_in) is
variable decimal: integer;
begin
decimal := to_integer(unsigned(data_in));
case(decimal) is
when 255 =>
x <= "00000010";
y <= "00000101";
n <="00000101";
when 254 =>
x <= "00000010";
y <= "00000101";
n <="00000100";
when 253 =>
x <= "00000010";
y <= "00000101";
n <="00000011";
when 252 =>
x <= "00000010";
y <= "00000101";
n <="00000010";
when 251 =>
x <= "00000010";
y <= "00000101";
n <="00000001";
when 250 =>
x <= "00000010";
y <= "00000101";
n <="00000000";
when 249 =>
x <= "00000010";
y <= "00000100";
n <="00001001";
when 248 =>
x <= "00000010";
y <= "00000100";
n <="00001000";
when 247 =>
x <= "00000010";
y <= "00000100";
n <="00000111";
when 246 =>
x <= "00000010";
y <= "00000100";
n <="00000110";
when 245 =>
x <= "00000010";
y <= "00000100";
n <="00000101";
when 244 =>
x <= "00000010";
y <= "00000100";
n <="00000100";
when 243 =>
x <= "00000010";
y <= "00000100";
n <="00000011";
when 242 =>
x <= "00000010";
y <= "00000100";
n <="00000010";
when 241 =>
x <= "00000010";
y <= "00000100";
n <="00000001";
when 240 =>
x <= "00000010";
y <= "00000100";
n <="00000000";
when 239 =>
x <= "00000010";
y <= "00000011";
n <="00001001";
when 238 =>
x <= "00000010";
y <= "00000011";
n <="00001000";
when 237 =>
x <= "00000010";
y <= "00000011";
n <="00000111";
when 236 =>
x <= "00000010";
y <= "00000011";
n <="00000110";
when 235 =>
x <= "00000010";
y <= "00000011";
n <="00000101";
when 234 =>
x <= "00000010";
y <= "00000011";
n <="00000100";
when 233 =>
x <= "00000010";
y <= "00000011";
n <="00000011";
when 232 =>
x <= "00000010";
y <= "00000011";
n <="00000010";
when 231 =>
x <= "00000010";
y <= "00000011";
n <="00000001";
when 230 =>
x <= "00000010";
y <= "00000011";
n <="00000000";
when 229 =>
x <= "00000010";
y <= "00000010";
n <="00001001";
when 228 =>
x <= "00000010";
y <= "00000010";
n <="00001000";
when 227 =>
x <= "00000010";
y <= "00000010";
n <="00000111";
when 226 =>
x <= "00000010";
y <= "00000010";
n <="00000110";
when 225 =>
x <= "00000010";
y <= "00000010";
n <="00000101";
when 224 =>
x <= "00000010";
y <= "00000010";
n <="00000100";
when 223 =>
x <= "00000010";
y <= "00000010";
n <="00000011";
when 222 =>
x <= "00000010";
y <= "00000010";
n <="00000010";
when 221 =>
x <= "00000010";
y <= "00000010";
n <="00000001";
when 220 =>
x <= "00000010";
y <= "00000010";
n <="00000000";
when 219 =>
x <= "00000010";
y <= "00000001";
n <="00001001";
when 218 =>
x <= "00000010";
y <= "00000001";
n <="00001000";
when 217 =>
x <= "00000010";
y <= "00000001";
n <="00000111";
when 216 =>
x <= "00000010";
y <= "00000001";
n <="00000110";
when 215 =>
x <= "00000010";
y <= "00000001";
n <="00000101";
when 214 =>
x <= "00000010";
y <= "00000001";
n <="00000100";
when 213 =>
x <= "00000010";
y <= "00000001";
n <="00000011";
when 212 =>
x <= "00000010";
y <= "00000001";
n <="00000010";
when 211 =>
x <= "00000010";
y <= "00000001";
n <="00000001";
when 210 =>
x <= "00000010";
y <= "00000001";
n <="00000000";
when 209 =>
x <= "00000010";
y <= "00000000";
n <="00001001";
when 208 =>
x <= "00000010";
y <= "00000000";
n <="00001000";
when 207 =>
x <= "00000010";
y <= "00000000";
n <="00000111";
when 206 =>
x <= "00000010";
y <= "00000000";
n <="00000110";
when 205 =>
x <= "00000010";
y <= "00000000";
n <="00000101";
when 204 =>
x <= "00000010";
y <= "00000000";
n <="00000100";
when 203 =>
x <= "00000010";
y <= "00000000";
n <="00000011";
when 202 =>
x <= "00000010";
y <= "00000000";
n <="00000010";
when 201 =>
x <= "00000010";
y <= "00000000";
n <="00000001";
when 200 =>
x <= "00000010";
y <= "00000000";
n <="00000000";
when 199 =>
x <= "00000001";
y <= "00001001";
n <="00001001";
when 198 =>
x <= "00000001";
y <= "00001001";
n <="00001000";
when 197 =>
x <= "00000001";
y <= "00001001";
n <="00000111";
when 196 =>
x <= "00000001";
y <= "00001001";
n <="00000110";
when 195 =>
x <= "00000001";
y <= "00001001";
n <="00000001";
when 194 =>
x <= "00000001";
y <= "00001001";
n <="00000100";
when 193 =>
x <= "00000001";
y <= "00001001";
n <="00000011";
when 192 =>
x <= "00000001";
y <= "00001001";
n <="00000010";
when 191 =>
x <= "00000001";
y <= "00001001";
n <="00000001";
when 190 =>
x <= "00000001";
y <= "00001001";
n <="00000000";
when 189 =>
x <= "00000001";
y <= "00001000";
n <="00001001";
when 188 =>
x <= "00000001";
y <= "00001000";
n <="00001000";
when 187 =>
x <= "00000001";
y <= "00001000";
n <="00000111";
when 186 =>
x <= "00000001";
y <= "00001000";
n <="00000110";
when 185 =>
x <= "00000001";
y <= "00001000";
n <="00000101";
when 184 =>
x <= "00000001";
y <= "00001000";
n <="00000100";
when 183 =>
x <= "00000001";
y <= "00001000";
n <="00000011";
when 182 =>
x <= "00000001";
y <= "00001000";
n <="00000010";
when 181 =>
x <= "00000001";
y <= "00001000";
n <= "00000001";
when 180 =>
x <= "00000001";
y <= "00001000";
n <="00000000";
when 179 =>
x <= "00000001";
y <= "00000111";
n <="00001001";
when 178 =>
x <= "00000001";
y <= "00000111";
n <="00001000";
when 177 =>
x <= "00000001";
y <= "00000111";
n <="00000111";
when 176 =>
x <= "00000001";
y <= "00000111";
n <="00000110";
when 175 =>
x <= "00000001";
y <= "00000111";
n <="00000101";
when 174 =>
x <= "00000001";
y <= "00000111";
n <="00000100";
when 173 =>
x <= "00000001";
y <= "00000111";
n <="00000011";
when 172 =>
x <= "00000001";
y <= "00000111";
n <="00000010";
when 171 =>
x <= "00000001";
y <= "00000111";
n <="00000001";
when 170 =>
x <= "00000001";
y <= "00000111";
n <="00000000";
when 169 =>
x <= "00000001";
y <= "00000110";
n <="00001001";
when 168 =>
x <= "00000001";
y <= "00000110";
n <="00001000";
when 167 =>
x <= "00000001";
y <= "00000110";
n <="00000111";
when 166 =>
x <= "00000001";
y <= "00000110";
n <="00000110";
when 165 =>
x <= "00000001";
y <= "00000110";
n <="00000101";
when 164 =>
x <= "00000001";
y <= "00000110";
n <="00000100";
when 163 =>
x <= "00000001";
y <= "00000110";
n <="00000011";
when 162 =>
x <= "00000001";
y <= "00000110";
n <="00000010";
when 161 =>
x <= "00000001";
y <= "00000110";
n <="00000001";
when 160 =>
x <= "00000001";
y <= "00000110";
n <="00000000";
when 159 =>
x <= "00000001";
y <= "00000101";
n <="00001001";
when 158 =>
x <= "00000001";
y <= "00000101";
n <="00001000";
when 157 =>
x <= "00000001";
y <= "00000101";
n <="00000111";
when 156 =>
x <= "00000001";
y <= "00000101";
n <="00000110";
when 155 =>
x <= "00000001";
y <= "00000101";
n <="00000101";
when 154 =>
x <= "00000001";
y <= "00000101";
n <="00000100";
when 153 =>
x <= "00000001";
y <= "00000101";
n <="00000011";
when 152 =>
x <= "00000001";
y <= "00000101";
n <="00000010";
when 151 =>
x <= "00000001";
y <= "00000101";
n <="00000001";
when 150 =>
x <= "00000001";
y <= "00000101";
n <="00000000";
when 149 =>
x <= "00000001";
y <= "00000100";
n <="00001001";
when 148 =>
x <= "00000001";
y <= "00000100";
n <="00001000";
when 147 =>
x <= "00000001";
y <= "00000100";
n <="00000111";
when 146 =>
x <= "00000001";
y <= "00000100";
n <="00000110";
when 145 =>
x <= "00000001";
y <= "00000100";
n <="00000101";
when 144 =>
x <= "00000001";
y <= "00000100";
n <="00000100";
when 143 =>
x <= "00000001";
y <= "00000100";
n <="00000011";
when 142 =>
x <= "00000001";
y <= "00000100";
n <="00000010";
when 141 =>
x <= "00000001";
y <= "00000100";
n <="00000001";
when 140 =>
x <= "00000001";
y <= "00000100";
n <="00000000";
when 139 =>
x <= "00000001";
y <= "00000011";
n <="00001001";
when 138 =>
x <= "00000001";
y <= "00000011";
n <="00001000";
when 137 =>
x <= "00000001";
y <= "00000011";
n <="00000111";
when 136 =>
x <= "00000001";
y <= "00000011";
n <="00000110";
when 135 =>
x <= "00000001";
y <= "00000011";
n <="00000101";
when 134 =>
x <= "00000001";
y <= "00000011";
n <="00000100";
when 133 =>
x <= "00000001";
y <= "00000011";
n <="00000101";
when 132 =>
x <= "00000001";
y <= "00000011";
n <="00000010";
when 131 =>
x <= "00000001";
y <= "00000011";
n <="00000001";
when 130 =>
x <= "00000001";
y <= "00000011";
n <="00000000";
when 129 =>
x <= "00000001";
y <= "00000010";
n <="00001001";
when 128 =>
x <= "00000001";
y <= "00000010";
n <="00001000";
when 127 =>
x <= "00000001";
y <= "00000010";
n <="00000111";
when 126 =>
x <= "00000001";
y <= "00000010";
n <="00000110";
when 125 =>
x <= "00000001";
y <= "00000010";
n <="00000101";
when 124 =>
x <= "00000001";
y <= "00000010";
n <="00000100";
when 123 =>
x <= "00000001";
y <= "00000010";
n <="00000011";
when 122 =>
x <= "00000001";
y <= "00000010";
n <="00000010";
when 121 =>
x <= "00000001";
y <= "00000010";
n <="00000001";
when 120 =>
x <= "00000001";
y <= "00000010";
n <="00000000";
when 119 =>
x <= "00000001";
y <= "00000001";
n <="00001001";
when 118 =>
x <= "00000001";
y <= "00000001";
n <="00001000";
when 117 =>
x <= "00000001";
y <= "00000001";
n <="00000111";
when 116 =>
x <= "00000001";
y <= "00000001";
n <="00000110";
when 115 =>
x <= "00000001";
y <= "00000001";
n <="00000101";
when 114 =>
x <= "00000001";
y <= "00000001";
n <="00000100";
when 113 =>
x <= "00000001";
y <= "00000001";
n <="00000011";
when 112 =>
x <= "00000001";
y <= "00000001";
n <="00000010";
when 111 =>
x <= "00000001";
y <= "00000001";
n <="00000001";
when 110 =>
x <= "00000001";
y <= "00000001";
n <="00000000";
when 109 =>
x <= "00000001";
y <= "00000000";
n <="00001001";
when 108 =>
x <= "00000001";
y <= "00000000";
n <="00001000";
when 107 =>
x <= "00000001";
y <= "00000000";
n <="00000111";
when 106 =>
x <= "00000001";
y <= "00000000";
n <="00000110";
when 105 =>
x <= "00000001";
y <= "00000000";
n <="00000101";
when 104 =>
x <= "00000001";
y <= "00000000";
n <="00000100";
when 103 =>
x <= "00000001";
y <= "00000000";
n <="00000011";
when 102 =>
x <= "00000001";
y <= "00000000";
n <="00000010";
when 101 =>
x <= "00000001";
y <= "00000000";
n <="00000001";
when 100 =>
x <= "00000001";
y <= "00000000";
n <="00000000";
when 99 =>
x <= "00000000";
y <= "00001001";
n <="00001001";
when 98 =>
x <= "00000000";
y <= "00001001";
n <="00001000";
when 97 =>
x <= "00000000";
y <= "00001001";
n <="00000111";
when 96 =>
x <= "00000000";
y <= "00001001";
n <="00000110";
when 95 =>
x <= "00000000";
y <= "00001001";
n <="00000101";
when 94 =>
x <= "00000000";
y <= "00001001";
n <="00000100";
when 93 =>
x <= "00000000";
y <= "00001001";
n <="00000011";
when 92 =>
x <= "00000000";
y <= "00001001";
n <="00000010";
when 91 =>
x <= "00000000";
y <= "00001001";
n <="00000001";
when 90 =>
x <= "00000000";
y <= "00001001";
n <="00000000";
when 89 =>
x <= "00000000";
y <= "00001000";
n <="00001001";
when 88 =>
x <= "00000000";
y <= "00001000";
n <="00001000";
when 87 =>
x <= "00000000";
y <= "00001000";
n <="00000111";
when 86 =>
x <= "00000000";
y <= "00001000";
n <="00000110";
when 85 =>
x <= "00000000";
y <= "00001000";
n <="00000100";
when 84 =>
x <= "00000000";
y <= "00001000";
n <="00000100";
when 83 =>
x <= "00000000";
y <= "00001000";
n <="00000011";
when 82 =>
x <= "00000000";
y <= "00001000";
n <="00000010";
when 81 =>
x <= "00000000";
y <= "00001000";
n <="00000001";
when 80 =>
x <= "00000000";
y <= "00001000";
n <="00000000";
when 79 =>
x <= "00000000";
y <= "00000111";
n <="00001001";
when 78 =>
x <= "00000000";
y <= "00000111";
n <="00001000";
when 77 =>
x <= "00000000";
y <= "00000111";
n <="00000111";
when 76 =>
x <= "00000000";
y <= "00000111";
n <="00000110";
when 75 =>
x <= "00000000";
y <= "00000111";
n <="00000101";
when 74 =>
x <= "00000000";
y <= "00000111";
n <="00000100";
when 73 =>
x <= "00000000";
y <= "00000111";
n <="00000011";
when 72 =>
x <= "00000000";
y <= "00000111";
n <="00000010";
when 71 =>
x <= "00000000";
y <= "00000111";
n <="00000001";
when 70 =>
x <= "00000000";
y <= "00000111";
n <="00000000";
when 69 =>
x <= "00000000";
y <= "00000110";
n <="00001001";
when 68 =>
x <= "00000000";
y <= "00000110";
n <="00001000";
when 67 =>
x <= "00000000";
y <= "00000110";
n <="00000111";
when 66 =>
x <= "00000000";
y <= "00000110";
n <="00000110";
when 65 =>
x <= "00000000";
y <= "00000110";
n <="00000101";
when 64 =>
x <= "00000000";
y <= "00000110";
n <="00000100";
when 63 =>
x <= "00000000";
y <= "00000110";
n <="00000011";
when 62 =>
x <= "00000000";
y <= "00000110";
n <="00000010";
when 61 =>
x <= "00000000";
y <= "00000110";
n <="00000001";
when 60 =>
x <= "00000000";
y <= "00000110";
n <="00000000";
when 59 =>
x <= "00000000";
y <= "00000101";
n <="00001001";
when 58 =>
x <= "00000000";
y <= "00000101";
n <="00001000";
when 57 =>
x <= "00000000";
y <= "00000101";
n <="00000111";
when 56 =>
x <= "00000000";
y <= "00000101";
n <="00000110";
when 55 =>
x <= "00000000";
y <= "00000101";
n <="00000101";
when 54 =>
x <= "00000000";
y <= "00000101";
n <="00000100";
when 53 =>
x <= "00000000";
y <= "00000101";
n <="00000011";
when 52 =>
x <= "00000000";
y <= "00000101";
n <="00000010";
when 51 =>
x <= "00000000";
y <= "00000101";
n <="00000001";
when 50 =>
x <= "00000000";
y <= "00000101";
n <="00000000";
when 49 =>
x <= "00000000";
y <= "00000100";
n <="00001001";
when 48 =>
x <= "00000000";
y <= "00000100";
n <="00001000";
when 47 =>
x <= "00000000";
y <= "00000100";
n <="00000111";
when 46 =>
x <= "00000000";
y <= "00000100";
n <="00000110";
when 45 =>
x <= "00000000";
y <= "00000100";
n <="00000101";
when 44 =>
x <= "00000000";
y <= "00000100";
n <="00000100";
when 43 =>
x <= "00000000";
y <= "00000100";
n <="00000011";
when 42 =>
x <= "00000000";
y <= "00000100";
n <="00000010";
when 41 =>
x <= "00000000";
y <= "00000100";
n <="00000001";
when 40 =>
x <= "00000000";
y <= "00000100";
n <="00000000";
when 39 =>
x <= "00000000";
y <= "00000011";
n <="00001001";
when 38 =>
x <= "00000000";
y <= "00000011";
n <="00001000";
when 37 =>
x <= "00000000";
y <= "00000011";
n <="00000111";
when 36 =>
x <= "00000000";
y <= "00000011";
n <="00000110";
when 35 =>
x <= "00000000";
y <= "00000011";
n <="00000101";
when 34 =>
x <= "00000000";
y <= "00000011";
n <="00000100";
when 33 =>
x <= "00000000";
y <= "00000011";
n <="00000011";
when 32 =>
x <= "00000000";
y <= "00000011";
n <="00000010";
when 31 =>
x <= "00000000";
y <= "00000011";
n <="00000001";
when 30 =>
x <= "00000000";
y <= "00000011";
n <="00000000";
when 29 =>
x <= "00000000";
y <= "00000010";
n <="00001001";
when 28 =>
x <= "00000000";
y <= "00000010";
n <="00001000";
when 27 =>
x <= "00000000";
y <= "00000010";
n <="00000111";
when 26 =>
x <= "00000000";
y <= "00000010";
n <="00000110";
when 25 =>
x <= "00000000";
y <= "00000010";
n <="00000000";
when 24 =>
x <= "00000000";
y <= "00000010";
n <="00000100";
when 23 =>
x <= "00000000";
y <= "00000010";
n <="00000011";
when 22 =>
x <= "00000000";
y <= "00000010";
n <="00000010";
when 21 =>
x <= "00000000";
y <= "00000010";
n <="00000001";
when 20 =>
x <= "00000000";
y <= "00000010";
n <="00000000";
when 19 =>
x <= "00000000";
y <= "00000001";
n <="00001001";
when 18 =>
x <= "00000000";
y <= "00000001";
n <="00001000";
when 17 =>
x <= "00000000";
y <= "00000001";
n <="00000111";
when 16 =>
x <= "00000000";
y <= "00000001";
n <="00000110";
when 15 =>
x <= "00000000";
y <= "00000001";
n <="00000101";
when 14 =>
x <= "00000000";
y <= "00000001";
n <="00000100";
when 13 =>
x <= "00000000";
y <= "00000001";
n <="00000011";
when 12 =>
x <= "00000000";
y <= "00000001";
n <="00000010";
when 11 =>
x <= "00000000";
y <= "00000001";
n <="00000001";
when 10 =>
x <= "00000000";
y <= "00000001";
n <="00000000";
when 9 =>
x <= "00000000";
y <= "00000000";
n <="00001001";
when 8 =>
x <= "00000000";
y <= "00000000";
n <="00001000";
when 7 =>
x <= "00000000";
y <= "00000000";
n <="00000111";
when 6 =>
x <= "00000000";
y <= "00000000";
n <="00000110";
when 5 =>
x <= "00000000";
y <= "00000000";
n <="00000101";
when 4 =>
x <= "00000000";
y <= "00000000";
n <="00000100";
when 3 =>
x <= "00000000";
y <= "00000000";
n <="00000011";
when 2 =>
x <= "00000000";
y <= "00000000";
n <="00000010";
when 1 =>
x <= "00000000";
y <= "00000000";
n <="00000001";
when 0 =>
x <= "00000000";
y <= "00000000";
n <="00000000";
when others =>
x <= "00000000";
y <= "00000000";
n <="00000000";
end case;
end process;

end Behavioral;
